`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

//
//////////////////////////////////////////////////////////////////////////////////
module mem256_16(clk, we, addr, d_in, d_out);
    

endmodule
